module clkbuffer(d_out,d_in);
input d_in;
output d_out;
buf(d_out,d_in);
endmodule